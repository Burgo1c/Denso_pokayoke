4,4,CODE39,M,16,IC04005512000001,1,,16,49433034303035353132303030303031,,,,,,�C�O�i�e�j
4,4,CODE39,M,10,IC04005512,1,,10,49433034303035353132,,,,,,�C�O�i�q�j
4,4,CODE39,M,16,6C05014510000001,1,,16,36433035303134353130303030303031,,,,,,�C�O�i�e�j
4,4,CODE39,M,10,6C05014510,1,,10,36433035303134353130,,,,,,�C�O�i�q�j
4,4,CODE39,M,16,1J55017322000001,1,,16,314A3535303137333232303030303031,,,,,,�C�O�i�e�j
4,4,CODE39,M,10,1J55017322,1,,10,314A3535303137333232,,,,,,�C�O�i�q�j
4,4,CODE39,M,10,PF80124950,1,,10,50463830313234393530,,,,,,����
4,4,CODE39,M,10,6C09054520,1,,10,36433039303534353230,,,,,,����
4,4,CODE39,M,10,3G74094202,1,,10,33473734303934323032,,,,,,����
